module control(
    input [6:0] ctrl,
    output branch,
    output RegWrite,
    output MemtoReg,
    output MemRead,
    output MemWrite,
    output alu_src,
    output [1:0] alu_op
);
    //alu op for 

endmodule