`include "alu.v"
`include "adder.v"
`include "alu_control.v"
`include "immgen.v"
`include "instruction_mem.v"
`include "control.v"
`include "mem.v"
`include "registers.v"

module (
    input clk; // clock control signal for the entire processor
);

// first, add the PC block connections



endmodule